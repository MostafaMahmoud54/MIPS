module And_Gate (
    input IN1,IN2,
    output wire AND_out
);

assign AND_out=IN1 & IN2;
endmodule